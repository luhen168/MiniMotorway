`timescale 1ns / 1ns
`define RVFI
import ibex_pkg::*;
module tb_ibex_riscv_compliance  #(
    // parameter bit          PMPEnable        = 1'b0,
    // parameter int unsigned PMPGranularity   = 0,
    // parameter int unsigned PMPNumRegions    = 4,
    // parameter int unsigned MHPMCounterNum   = 0,
    // parameter int unsigned MHPMCounterWidth = 40,
    // parameter bit RV32E                     = 1'b0,
    // parameter ibex_pkg::rv32m_e RV32M       = ibex_pkg::RV32MNone,
    // parameter ibex_pkg::rv32b_e RV32B       = ibex_pkg::RV32BNone,
    // parameter ibex_pkg::regfile_e RegFile   = ibex_pkg::RegFileFF,
    // parameter bit BranchTargetALU           = 1'b0,
    // parameter bit WritebackStage            = 1'b0,
    // parameter bit ICache                    = 1'b0,
    // parameter bit ICacheECC                 = 1'b0,
    // parameter bit BranchPredictor           = 1'b0,
    // parameter bit SecureIbex                = 1'b0,
    // parameter bit ICacheScramble            = 1'b0,
    // parameter bit DbgTriggerEn              = 1'b0
) (
  
);

    logic clk_sys_i, rst_sys_ni;

      // Instantiate the ibex_top
  ibex_riscv_compliance u_ibex_riscv_compliance_i(
      .IO_CLK(clk_sys_i),
      .IO_RST_N(rst_sys_ni)
  );

  // Clock generation
  initial begin
    clk_sys_i = 0;
    forever #5 clk_sys_i = ~clk_sys_i;
  end

  // Test sequence
  initial begin
    // Initialize inputs
    rst_sys_ni = 0;
    // Release reset after some time
    #10 rst_sys_ni = 1;
    //Stop simulation
    repeat (100000) @(posedge clk_sys_i);
    $stop;
  end

endmodule 