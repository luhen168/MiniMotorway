module if_stage #(
    parameters
) (
    // Signal synchronous (clk) and acsynchronous (rst)
    input clk,
    input rst,

    // 


);
    
endmodule